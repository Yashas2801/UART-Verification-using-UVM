module top;
  import uvm_pkg::*;
  import UART_pkg::*;

  initial begin
    run_test();
  end
endmodule
