`timescale 1ns / 10ps
package UART_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "xtn.sv"
  `include "agent_config.sv"
  `include "env_config.sv"
  `include "sequence.sv"

  `include "driver.sv"
  `include "monitor.sv"
  `include "sequencer.sv"
  `include "agent.sv"

  `include "virtual_sequencer.sv"
  `include "virtual_sequence.sv"

  `include "env.sv"
  `include "test.sv"

endpackage
